module traffic_system_top (
    input clk,
    input rst_n,
    input traffic_jam_0;
    input traffic_jam_1;
    input traffic_jam_2;
    input traffic_jam_3;
    output reg allow_0;
    output reg allow_1;
    output reg allow_2;
    output reg allow_3;
);
    
endmodule